   
    parameter PROC_NUM = 52;
    parameter ST_IDLE = 3'b000;
    parameter ST_FILTER_FAKE = 3'b001;
    parameter ST_DL_DETECTED = 3'b010;
    parameter ST_DL_REPORT = 3'b100;
   

    reg [2:0] CS_fsm;
    reg [2:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    reg [31:0] dl_keep_cnt;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg or dl_keep_cnt) begin
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_FILTER_FAKE;
                end
                else begin
                    NS_fsm = ST_IDLE;
                end
            end
            ST_FILTER_FAKE: begin
                if (dl_keep_cnt >= 32'd1000) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else if (dl_detect_reg != (dl_detect_reg & dl_in_vec)) begin
                    NS_fsm = ST_IDLE;
                end
                else begin
                    NS_fsm = ST_FILTER_FAKE;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
                else begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            default: NS_fsm = ST_IDLE;
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_keep_cnt <= 32'h0;
        end
        else begin
            if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg == (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= dl_keep_cnt + 32'h1;
            end
            else if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg != (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= 32'h0;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = (|dl_detect_reg) && (CS_fsm == ST_DL_DETECTED || CS_fsm == ST_DL_REPORT);

    // dl_done_reg record the cycles has been reported
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    wire [PROC_NUM*PROC_NUM - 1:0] origin_tmp;
    assign origin_tmp[PROC_NUM - 1:0] = (dl_detect_reg[0] & ~dl_done_reg[0]) ? 'b1 : 'b0;
    genvar j;
    generate
    for(j = 1;j < PROC_NUM;j = j + 1) begin: F1
        assign origin_tmp[j*PROC_NUM +: PROC_NUM] = (dl_detect_reg[j] & ~dl_done_reg[j]) ? ('b1 << j) : origin_tmp[(j - 1)*PROC_NUM +: PROC_NUM];
    end
    endgenerate
    always @ (CS_fsm or origin_tmp) begin
        if (CS_fsm == ST_DL_DETECTED) begin
            origin = origin_tmp[(PROC_NUM - 1)*PROC_NUM +: PROC_NUM];
        end
        else begin
            origin = 'b0;
        end
    end

    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // find_df_deadlock to report the deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            find_df_deadlock <= 1'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED && dl_detect_reg == dl_done_reg) begin
                find_df_deadlock <= 1'b1;
            end
            else if (CS_fsm == ST_IDLE) begin
                find_df_deadlock <= 1'b0;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [560:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "rocev2_top_rocev2_top.entry_proc_U0";
                end
                1 : begin
                    proc_path = "rocev2_top_rocev2_top.convert_axis_to_net_axis_512_U0";
                end
                2 : begin
                    proc_path = "rocev2_top_rocev2_top.convert_net_axis_to_axis_512_U0";
                end
                3 : begin
                    proc_path = "rocev2_top_rocev2_top.convert_axis_to_net_axis_512_1_U0";
                end
                4 : begin
                    proc_path = "rocev2_top_rocev2_top.convert_net_axis_to_axis_512_2_U0";
                end
                5 : begin
                    proc_path = "rocev2_top_rocev2_top.extract_icrc_512_0_U0";
                end
                6 : begin
                    proc_path = "rocev2_top_rocev2_top.insert_icrc_512_0_U0";
                end
                7 : begin
                    proc_path = "rocev2_top_rocev2_top.process_ipv4_512_U0";
                end
                8 : begin
                    proc_path = "rocev2_top_rocev2_top.ipv4_drop_optional_ip_header_512_U0";
                end
                9 : begin
                    proc_path = "rocev2_top_rocev2_top.ipv4_lshiftWordByOctet_512_2_U0";
                end
                10 : begin
                    proc_path = "rocev2_top_rocev2_top.ipv4_generate_ipv4_512_3_U0";
                end
                11 : begin
                    proc_path = "rocev2_top_rocev2_top.process_udp_512_4_U0";
                end
                12 : begin
                    proc_path = "rocev2_top_rocev2_top.udp_rshiftWordByOctet_net_axis_512_512_2_U0";
                end
                13 : begin
                    proc_path = "rocev2_top_rocev2_top.merge_rx_meta_U0";
                end
                14 : begin
                    proc_path = "rocev2_top_rocev2_top.split_tx_meta_U0";
                end
                15 : begin
                    proc_path = "rocev2_top_rocev2_top.udp_lshiftWordByOctet_512_1_U0";
                end
                16 : begin
                    proc_path = "rocev2_top_rocev2_top.generate_udp_512_U0";
                end
                17 : begin
                    proc_path = "rocev2_top_rocev2_top.qp_interface_0_U0";
                end
                18 : begin
                    proc_path = "rocev2_top_rocev2_top.rx_process_ibh_512_0_U0";
                end
                19 : begin
                    proc_path = "rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_11_0_U0";
                end
                20 : begin
                    proc_path = "rocev2_top_rocev2_top.rx_process_exh_512_0_U0";
                end
                21 : begin
                    proc_path = "rocev2_top_rocev2_top.rx_ibh_fsm_0_U0";
                end
                22 : begin
                    proc_path = "rocev2_top_rocev2_top.drop_ooo_ibh_512_0_U0";
                end
                23 : begin
                    proc_path = "rocev2_top_rocev2_top.ipUdpMetaHandler_512_0_U0";
                end
                24 : begin
                    proc_path = "rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0";
                end
                25 : begin
                    proc_path = "rocev2_top_rocev2_top.rx_exh_payload_512_0_U0";
                end
                26 : begin
                    proc_path = "rocev2_top_rocev2_top.handle_read_requests_0_U0";
                end
                27 : begin
                    proc_path = "rocev2_top_rocev2_top.stream_merger_ackEvent_U0";
                end
                28 : begin
                    proc_path = "rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_12_0_U0";
                end
                29 : begin
                    proc_path = "rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_13_0_U0";
                end
                30 : begin
                    proc_path = "rocev2_top_rocev2_top.merge_rx_pkgs_512_0_U0";
                end
                31 : begin
                    proc_path = "rocev2_top_rocev2_top.local_req_handler_0_U0";
                end
                32 : begin
                    proc_path = "rocev2_top_rocev2_top.tx_pkg_arbiter_512_0_U0";
                end
                33 : begin
                    proc_path = "rocev2_top_rocev2_top.meta_merger_0_U0";
                end
                34 : begin
                    proc_path = "rocev2_top_rocev2_top.lshiftWordByOctet_512_12_0_U0";
                end
                35 : begin
                    proc_path = "rocev2_top_rocev2_top.lshiftWordByOctet_512_13_0_U0";
                end
                36 : begin
                    proc_path = "rocev2_top_rocev2_top.generate_exh_512_0_U0";
                end
                37 : begin
                    proc_path = "rocev2_top_rocev2_top.append_payload_512_0_U0";
                end
                38 : begin
                    proc_path = "rocev2_top_rocev2_top.lshiftWordByOctet_512_11_0_U0";
                end
                39 : begin
                    proc_path = "rocev2_top_rocev2_top.generate_ibh_512_0_U0";
                end
                40 : begin
                    proc_path = "rocev2_top_rocev2_top.prepend_ibh_header_512_0_U0";
                end
                41 : begin
                    proc_path = "rocev2_top_rocev2_top.tx_ipUdpMetaMerger_0_U0";
                end
                42 : begin
                    proc_path = "rocev2_top_rocev2_top.mem_cmd_merger_512_0_U0";
                end
                43 : begin
                    proc_path = "rocev2_top_rocev2_top.conn_table_0_U0";
                end
                44 : begin
                    proc_path = "rocev2_top_rocev2_top.state_table_0_U0";
                end
                45 : begin
                    proc_path = "rocev2_top_rocev2_top.msn_table_0_U0";
                end
                46 : begin
                    proc_path = "rocev2_top_rocev2_top.merge_retrans_request_U0";
                end
                47 : begin
                    proc_path = "rocev2_top_rocev2_top.transport_timer_0_U0";
                end
                48 : begin
                    proc_path = "rocev2_top_rocev2_top.freelist_handler_0_U0";
                end
                49 : begin
                    proc_path = "rocev2_top_rocev2_top.retrans_pointer_table_0_U0";
                end
                50 : begin
                    proc_path = "rocev2_top_rocev2_top.retrans_meta_table_0_U0";
                end
                51 : begin
                    proc_path = "rocev2_top_rocev2_top.process_retransmissions_0_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [560:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num, input integer record_time);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", record_time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [560:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [472:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    10: begin
                        if (~entry_proc_U0.local_ip_address_c_blk_n) begin
                            if (~local_ip_address_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.local_ip_address_c_U' written by process 'rocev2_top_rocev2_top.ipv4_generate_ipv4_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.local_ip_address_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~local_ip_address_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.local_ip_address_c_U' read by process 'rocev2_top_rocev2_top.ipv4_generate_ipv4_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.local_ip_address_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    5: begin
                        if (~convert_axis_to_net_axis_512_U0.s_axis_rx_data_internal_blk_n) begin
                            if (~s_axis_rx_data_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.s_axis_rx_data_internal_U' written by process 'rocev2_top_rocev2_top.extract_icrc_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.s_axis_rx_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~s_axis_rx_data_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.s_axis_rx_data_internal_U' read by process 'rocev2_top_rocev2_top.extract_icrc_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.s_axis_rx_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                2 : begin
                    case(index2)
                    6: begin
                        if (~convert_net_axis_to_axis_512_U0.m_axis_tx_data_internal_blk_n) begin
                            if (~m_axis_tx_data_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.m_axis_tx_data_internal_U' written by process 'rocev2_top_rocev2_top.insert_icrc_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.m_axis_tx_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~m_axis_tx_data_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.m_axis_tx_data_internal_U' read by process 'rocev2_top_rocev2_top.insert_icrc_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.m_axis_tx_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                3 : begin
                    case(index2)
                    32: begin
                        if (~convert_axis_to_net_axis_512_1_U0.s_axis_mem_read_data_internal_blk_n) begin
                            if (~s_axis_mem_read_data_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.s_axis_mem_read_data_internal_U' written by process 'rocev2_top_rocev2_top.tx_pkg_arbiter_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.s_axis_mem_read_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~s_axis_mem_read_data_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.s_axis_mem_read_data_internal_U' read by process 'rocev2_top_rocev2_top.tx_pkg_arbiter_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.s_axis_mem_read_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                4 : begin
                    case(index2)
                    30: begin
                        if (~convert_net_axis_to_axis_512_2_U0.m_axis_mem_write_data_internal_blk_n) begin
                            if (~m_axis_mem_write_data_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.m_axis_mem_write_data_internal_U' written by process 'rocev2_top_rocev2_top.merge_rx_pkgs_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.m_axis_mem_write_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~m_axis_mem_write_data_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.m_axis_mem_write_data_internal_U' read by process 'rocev2_top_rocev2_top.merge_rx_pkgs_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.m_axis_mem_write_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                5 : begin
                    case(index2)
                    1: begin
                        if (~extract_icrc_512_0_U0.s_axis_rx_data_internal_blk_n) begin
                            if (~s_axis_rx_data_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.s_axis_rx_data_internal_U' written by process 'rocev2_top_rocev2_top.convert_axis_to_net_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.s_axis_rx_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~s_axis_rx_data_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.s_axis_rx_data_internal_U' read by process 'rocev2_top_rocev2_top.convert_axis_to_net_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.s_axis_rx_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    7: begin
                        if (~extract_icrc_512_0_U0.rx_crc2ipFifo_blk_n) begin
                            if (~rx_crc2ipFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_crc2ipFifo_U' written by process 'rocev2_top_rocev2_top.process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_crc2ipFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_crc2ipFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_crc2ipFifo_U' read by process 'rocev2_top_rocev2_top.process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_crc2ipFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                6 : begin
                    case(index2)
                    10: begin
                        if (~insert_icrc_512_0_U0.tx_ip2crcFifo_blk_n) begin
                            if (~tx_ip2crcFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_ip2crcFifo_U' written by process 'rocev2_top_rocev2_top.ipv4_generate_ipv4_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ip2crcFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_ip2crcFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_ip2crcFifo_U' read by process 'rocev2_top_rocev2_top.ipv4_generate_ipv4_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ip2crcFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (~insert_icrc_512_0_U0.m_axis_tx_data_internal_blk_n) begin
                            if (~m_axis_tx_data_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.m_axis_tx_data_internal_U' written by process 'rocev2_top_rocev2_top.convert_net_axis_to_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.m_axis_tx_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~m_axis_tx_data_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.m_axis_tx_data_internal_U' read by process 'rocev2_top_rocev2_top.convert_net_axis_to_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.m_axis_tx_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                7 : begin
                    case(index2)
                    5: begin
                        if (~process_ipv4_512_U0.rx_crc2ipFifo_blk_n) begin
                            if (~rx_crc2ipFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_crc2ipFifo_U' written by process 'rocev2_top_rocev2_top.extract_icrc_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_crc2ipFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_crc2ipFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_crc2ipFifo_U' read by process 'rocev2_top_rocev2_top.extract_icrc_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_crc2ipFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    8: begin
                        if (~process_ipv4_512_U0.rx_process2dropFifo_blk_n) begin
                            if (~rx_process2dropFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_process2dropFifo_U' written by process 'rocev2_top_rocev2_top.ipv4_drop_optional_ip_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_process2dropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_process2dropFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_process2dropFifo_U' read by process 'rocev2_top_rocev2_top.ipv4_drop_optional_ip_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_process2dropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~process_ipv4_512_U0.rx_process2dropLengthFifo_blk_n) begin
                            if (~rx_process2dropLengthFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_process2dropLengthFifo_U' written by process 'rocev2_top_rocev2_top.ipv4_drop_optional_ip_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_process2dropLengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_process2dropLengthFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_process2dropLengthFifo_U' read by process 'rocev2_top_rocev2_top.ipv4_drop_optional_ip_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_process2dropLengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~process_ipv4_512_U0.rx_ip2udpMetaFifo_blk_n) begin
                            if (~rx_ip2udpMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ip2udpMetaFifo_U' written by process 'rocev2_top_rocev2_top.merge_rx_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ip2udpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ip2udpMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ip2udpMetaFifo_U' read by process 'rocev2_top_rocev2_top.merge_rx_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ip2udpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                8 : begin
                    case(index2)
                    7: begin
                        if (~ipv4_drop_optional_ip_header_512_U0.rx_process2dropLengthFifo_blk_n) begin
                            if (~rx_process2dropLengthFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_process2dropLengthFifo_U' written by process 'rocev2_top_rocev2_top.process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_process2dropLengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_process2dropLengthFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_process2dropLengthFifo_U' read by process 'rocev2_top_rocev2_top.process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_process2dropLengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~ipv4_drop_optional_ip_header_512_U0.rx_process2dropFifo_blk_n) begin
                            if (~rx_process2dropFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_process2dropFifo_U' written by process 'rocev2_top_rocev2_top.process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_process2dropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_process2dropFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_process2dropFifo_U' read by process 'rocev2_top_rocev2_top.process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_process2dropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    11: begin
                        if (~ipv4_drop_optional_ip_header_512_U0.rx_ip2udpFifo_blk_n) begin
                            if (~rx_ip2udpFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ip2udpFifo_U' written by process 'rocev2_top_rocev2_top.process_udp_512_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ip2udpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ip2udpFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ip2udpFifo_U' read by process 'rocev2_top_rocev2_top.process_udp_512_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ip2udpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                9 : begin
                    case(index2)
                    10: begin
                        if (~ipv4_lshiftWordByOctet_512_2_U0.tx_shift2ipv4Fifo_blk_n) begin
                            if (~tx_shift2ipv4Fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_shift2ipv4Fifo_U' written by process 'rocev2_top_rocev2_top.ipv4_generate_ipv4_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_shift2ipv4Fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_shift2ipv4Fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_shift2ipv4Fifo_U' read by process 'rocev2_top_rocev2_top.ipv4_generate_ipv4_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_shift2ipv4Fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    16: begin
                        if (~ipv4_lshiftWordByOctet_512_2_U0.tx_udp2ipFifo_blk_n) begin
                            if (~tx_udp2ipFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_udp2ipFifo_U' written by process 'rocev2_top_rocev2_top.generate_udp_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_udp2ipFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_udp2ipFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_udp2ipFifo_U' read by process 'rocev2_top_rocev2_top.generate_udp_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_udp2ipFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                10 : begin
                    case(index2)
                    0: begin
                        if (~ipv4_generate_ipv4_512_3_U0.local_ip_address_blk_n) begin
                            if (~local_ip_address_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.local_ip_address_c_U' written by process 'rocev2_top_rocev2_top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.local_ip_address_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~local_ip_address_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.local_ip_address_c_U' read by process 'rocev2_top_rocev2_top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.local_ip_address_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (~ipv4_generate_ipv4_512_3_U0.tx_udp2ipMetaFifo_blk_n) begin
                            if (~tx_udp2ipMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_udp2ipMetaFifo_U' written by process 'rocev2_top_rocev2_top.split_tx_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_udp2ipMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_udp2ipMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_udp2ipMetaFifo_U' read by process 'rocev2_top_rocev2_top.split_tx_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_udp2ipMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    6: begin
                        if (~ipv4_generate_ipv4_512_3_U0.tx_ip2crcFifo_blk_n) begin
                            if (~tx_ip2crcFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_ip2crcFifo_U' written by process 'rocev2_top_rocev2_top.insert_icrc_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ip2crcFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_ip2crcFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_ip2crcFifo_U' read by process 'rocev2_top_rocev2_top.insert_icrc_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ip2crcFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    9: begin
                        if (~ipv4_generate_ipv4_512_3_U0.tx_shift2ipv4Fifo_blk_n) begin
                            if (~tx_shift2ipv4Fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_shift2ipv4Fifo_U' written by process 'rocev2_top_rocev2_top.ipv4_lshiftWordByOctet_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_shift2ipv4Fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_shift2ipv4Fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_shift2ipv4Fifo_U' read by process 'rocev2_top_rocev2_top.ipv4_lshiftWordByOctet_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_shift2ipv4Fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                11 : begin
                    case(index2)
                    8: begin
                        if (~process_udp_512_4_U0.rx_ip2udpFifo_blk_n) begin
                            if (~rx_ip2udpFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ip2udpFifo_U' written by process 'rocev2_top_rocev2_top.ipv4_drop_optional_ip_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ip2udpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ip2udpFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ip2udpFifo_U' read by process 'rocev2_top_rocev2_top.ipv4_drop_optional_ip_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ip2udpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    12: begin
                        if (~process_udp_512_4_U0.rx_udp2shiftFifo_blk_n) begin
                            if (~rx_udp2shiftFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_udp2shiftFifo_U' written by process 'rocev2_top_rocev2_top.udp_rshiftWordByOctet_net_axis_512_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_udp2shiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_udp2shiftFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_udp2shiftFifo_U' read by process 'rocev2_top_rocev2_top.udp_rshiftWordByOctet_net_axis_512_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_udp2shiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~process_udp_512_4_U0.rx_udpMetaFifo_blk_n) begin
                            if (~rx_udpMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_udpMetaFifo_U' written by process 'rocev2_top_rocev2_top.merge_rx_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_udpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_udpMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_udpMetaFifo_U' read by process 'rocev2_top_rocev2_top.merge_rx_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_udpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                12 : begin
                    case(index2)
                    11: begin
                        if (~udp_rshiftWordByOctet_net_axis_512_512_2_U0.rx_udp2shiftFifo_blk_n) begin
                            if (~rx_udp2shiftFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_udp2shiftFifo_U' written by process 'rocev2_top_rocev2_top.process_udp_512_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_udp2shiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_udp2shiftFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_udp2shiftFifo_U' read by process 'rocev2_top_rocev2_top.process_udp_512_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_udp2shiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    18: begin
                        if (~udp_rshiftWordByOctet_net_axis_512_512_2_U0.rx_udp2ibFifo_blk_n) begin
                            if (~rx_udp2ibFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_udp2ibFifo_U' written by process 'rocev2_top_rocev2_top.rx_process_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_udp2ibFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_udp2ibFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_udp2ibFifo_U' read by process 'rocev2_top_rocev2_top.rx_process_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_udp2ibFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                13 : begin
                    case(index2)
                    7: begin
                        if (~merge_rx_meta_U0.rx_ip2udpMetaFifo_blk_n) begin
                            if (~rx_ip2udpMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ip2udpMetaFifo_U' written by process 'rocev2_top_rocev2_top.process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ip2udpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ip2udpMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ip2udpMetaFifo_U' read by process 'rocev2_top_rocev2_top.process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ip2udpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    11: begin
                        if (~merge_rx_meta_U0.rx_udpMetaFifo_blk_n) begin
                            if (~rx_udpMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_udpMetaFifo_U' written by process 'rocev2_top_rocev2_top.process_udp_512_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_udpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_udpMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_udpMetaFifo_U' read by process 'rocev2_top_rocev2_top.process_udp_512_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_udpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    23: begin
                        if (~merge_rx_meta_U0.rx_ipUdpMetaFifo_blk_n) begin
                            if (~rx_ipUdpMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ipUdpMetaFifo_U' written by process 'rocev2_top_rocev2_top.ipUdpMetaHandler_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ipUdpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ipUdpMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ipUdpMetaFifo_U' read by process 'rocev2_top_rocev2_top.ipUdpMetaHandler_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ipUdpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                14 : begin
                    case(index2)
                    41: begin
                        if (~split_tx_meta_U0.tx_ipUdpMetaFifo_blk_n) begin
                            if (~tx_ipUdpMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_ipUdpMetaFifo_U' written by process 'rocev2_top_rocev2_top.tx_ipUdpMetaMerger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ipUdpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_ipUdpMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_ipUdpMetaFifo_U' read by process 'rocev2_top_rocev2_top.tx_ipUdpMetaMerger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ipUdpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    10: begin
                        if (~split_tx_meta_U0.tx_udp2ipMetaFifo_blk_n) begin
                            if (~tx_udp2ipMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_udp2ipMetaFifo_U' written by process 'rocev2_top_rocev2_top.ipv4_generate_ipv4_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_udp2ipMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_udp2ipMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_udp2ipMetaFifo_U' read by process 'rocev2_top_rocev2_top.ipv4_generate_ipv4_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_udp2ipMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    16: begin
                        if (~split_tx_meta_U0.tx_udpMetaFifo_blk_n) begin
                            if (~tx_udpMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_udpMetaFifo_U' written by process 'rocev2_top_rocev2_top.generate_udp_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_udpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_udpMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_udpMetaFifo_U' read by process 'rocev2_top_rocev2_top.generate_udp_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_udpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                15 : begin
                    case(index2)
                    16: begin
                        if (~udp_lshiftWordByOctet_512_1_U0.tx_shift2udpFifo_blk_n) begin
                            if (~tx_shift2udpFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_shift2udpFifo_U' written by process 'rocev2_top_rocev2_top.generate_udp_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_shift2udpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_shift2udpFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_shift2udpFifo_U' read by process 'rocev2_top_rocev2_top.generate_udp_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_shift2udpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    40: begin
                        if (~udp_lshiftWordByOctet_512_1_U0.tx_ib2udpFifo_blk_n) begin
                            if (~tx_ib2udpFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_ib2udpFifo_U' written by process 'rocev2_top_rocev2_top.prepend_ibh_header_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ib2udpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_ib2udpFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_ib2udpFifo_U' read by process 'rocev2_top_rocev2_top.prepend_ibh_header_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ib2udpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                16 : begin
                    case(index2)
                    14: begin
                        if (~generate_udp_512_U0.tx_udpMetaFifo_blk_n) begin
                            if (~tx_udpMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_udpMetaFifo_U' written by process 'rocev2_top_rocev2_top.split_tx_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_udpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_udpMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_udpMetaFifo_U' read by process 'rocev2_top_rocev2_top.split_tx_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_udpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    9: begin
                        if (~generate_udp_512_U0.tx_udp2ipFifo_blk_n) begin
                            if (~tx_udp2ipFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_udp2ipFifo_U' written by process 'rocev2_top_rocev2_top.ipv4_lshiftWordByOctet_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_udp2ipFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_udp2ipFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_udp2ipFifo_U' read by process 'rocev2_top_rocev2_top.ipv4_lshiftWordByOctet_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_udp2ipFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    15: begin
                        if (~generate_udp_512_U0.tx_shift2udpFifo_blk_n) begin
                            if (~tx_shift2udpFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_shift2udpFifo_U' written by process 'rocev2_top_rocev2_top.udp_lshiftWordByOctet_512_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_shift2udpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_shift2udpFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_shift2udpFifo_U' read by process 'rocev2_top_rocev2_top.udp_lshiftWordByOctet_512_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_shift2udpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                17 : begin
                    case(index2)
                    44: begin
                        if (~qp_interface_0_U0.qpi2stateTable_upd_req_blk_n) begin
                            if (~qpi2stateTable_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.qpi2stateTable_upd_req_U' written by process 'rocev2_top_rocev2_top.state_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.qpi2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~qpi2stateTable_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.qpi2stateTable_upd_req_U' read by process 'rocev2_top_rocev2_top.state_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.qpi2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~qp_interface_0_U0.stateTable2qpi_rsp_blk_n) begin
                            if (~stateTable2qpi_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.stateTable2qpi_rsp_U' written by process 'rocev2_top_rocev2_top.state_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.stateTable2qpi_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2qpi_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.stateTable2qpi_rsp_U' read by process 'rocev2_top_rocev2_top.state_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.stateTable2qpi_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    45: begin
                        if (~qp_interface_0_U0.if2msnTable_init_blk_n) begin
                            if (~if2msnTable_init_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.if2msnTable_init_U' written by process 'rocev2_top_rocev2_top.msn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.if2msnTable_init_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~if2msnTable_init_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.if2msnTable_init_U' read by process 'rocev2_top_rocev2_top.msn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.if2msnTable_init_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                18 : begin
                    case(index2)
                    12: begin
                        if (~rx_process_ibh_512_0_U0.rx_udp2ibFifo_blk_n) begin
                            if (~rx_udp2ibFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_udp2ibFifo_U' written by process 'rocev2_top_rocev2_top.udp_rshiftWordByOctet_net_axis_512_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_udp2ibFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_udp2ibFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_udp2ibFifo_U' read by process 'rocev2_top_rocev2_top.udp_rshiftWordByOctet_net_axis_512_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_udp2ibFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (~rx_process_ibh_512_0_U0.rx_ibh2shiftFifo_blk_n) begin
                            if (~rx_ibh2shiftFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibh2shiftFifo_U' written by process 'rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_11_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibh2shiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibh2shiftFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibh2shiftFifo_U' read by process 'rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_11_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibh2shiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    21: begin
                        if (~rx_process_ibh_512_0_U0.rx_ibh2fsm_MetaFifo_blk_n) begin
                            if (~rx_ibh2fsm_MetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibh2fsm_MetaFifo_U' written by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibh2fsm_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibh2fsm_MetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibh2fsm_MetaFifo_U' read by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibh2fsm_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (~rx_process_ibh_512_0_U0.rx_ibh2exh_MetaFifo_blk_n) begin
                            if (~rx_ibh2exh_MetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibh2exh_MetaFifo_U' written by process 'rocev2_top_rocev2_top.rx_process_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibh2exh_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibh2exh_MetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibh2exh_MetaFifo_U' read by process 'rocev2_top_rocev2_top.rx_process_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibh2exh_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                19 : begin
                    case(index2)
                    18: begin
                        if (~rshiftWordByOctet_net_axis_512_512_11_0_U0.rx_ibh2shiftFifo_blk_n) begin
                            if (~rx_ibh2shiftFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibh2shiftFifo_U' written by process 'rocev2_top_rocev2_top.rx_process_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibh2shiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibh2shiftFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibh2shiftFifo_U' read by process 'rocev2_top_rocev2_top.rx_process_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibh2shiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (~rshiftWordByOctet_net_axis_512_512_11_0_U0.rx_shift2exhFifo_blk_n) begin
                            if (~rx_shift2exhFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_shift2exhFifo_U' written by process 'rocev2_top_rocev2_top.rx_process_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_shift2exhFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_shift2exhFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_shift2exhFifo_U' read by process 'rocev2_top_rocev2_top.rx_process_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_shift2exhFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                20 : begin
                    case(index2)
                    18: begin
                        if (~rx_process_exh_512_0_U0.rx_ibh2exh_MetaFifo_blk_n) begin
                            if (~rx_ibh2exh_MetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibh2exh_MetaFifo_U' written by process 'rocev2_top_rocev2_top.rx_process_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibh2exh_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibh2exh_MetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibh2exh_MetaFifo_U' read by process 'rocev2_top_rocev2_top.rx_process_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibh2exh_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (~rx_process_exh_512_0_U0.rx_shift2exhFifo_blk_n) begin
                            if (~rx_shift2exhFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_shift2exhFifo_U' written by process 'rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_11_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_shift2exhFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_shift2exhFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_shift2exhFifo_U' read by process 'rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_11_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_shift2exhFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    22: begin
                        if (~rx_process_exh_512_0_U0.rx_exh2dropFifo_blk_n) begin
                            if (~rx_exh2dropFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exh2dropFifo_U' written by process 'rocev2_top_rocev2_top.drop_ooo_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2dropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exh2dropFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exh2dropFifo_U' read by process 'rocev2_top_rocev2_top.drop_ooo_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2dropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    21: begin
                        if (~rx_process_exh_512_0_U0.rx_exhMetaFifo_blk_n) begin
                            if (~rx_exhMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exhMetaFifo_U' written by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exhMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exhMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exhMetaFifo_U' read by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exhMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    23: begin
                        if (~rx_process_exh_512_0_U0.rx_exh2drop_MetaFifo_blk_n) begin
                            if (~rx_exh2drop_MetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exh2drop_MetaFifo_U' written by process 'rocev2_top_rocev2_top.ipUdpMetaHandler_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2drop_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exh2drop_MetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exh2drop_MetaFifo_U' read by process 'rocev2_top_rocev2_top.ipUdpMetaHandler_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2drop_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                21 : begin
                    case(index2)
                    18: begin
                        if (~rx_ibh_fsm_0_U0.rx_ibh2fsm_MetaFifo_blk_n) begin
                            if (~rx_ibh2fsm_MetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibh2fsm_MetaFifo_U' written by process 'rocev2_top_rocev2_top.rx_process_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibh2fsm_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibh2fsm_MetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibh2fsm_MetaFifo_U' read by process 'rocev2_top_rocev2_top.rx_process_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibh2fsm_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (~rx_ibh_fsm_0_U0.rx_exhMetaFifo_blk_n) begin
                            if (~rx_exhMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exhMetaFifo_U' written by process 'rocev2_top_rocev2_top.rx_process_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exhMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exhMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exhMetaFifo_U' read by process 'rocev2_top_rocev2_top.rx_process_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exhMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    44: begin
                        if (~rx_ibh_fsm_0_U0.rxIbh2stateTable_upd_req_blk_n) begin
                            if (~rxIbh2stateTable_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rxIbh2stateTable_upd_req_U' written by process 'rocev2_top_rocev2_top.state_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rxIbh2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxIbh2stateTable_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rxIbh2stateTable_upd_req_U' read by process 'rocev2_top_rocev2_top.state_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rxIbh2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rx_ibh_fsm_0_U0.stateTable2rxIbh_rsp_blk_n) begin
                            if (~stateTable2rxIbh_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.stateTable2rxIbh_rsp_U' written by process 'rocev2_top_rocev2_top.state_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.stateTable2rxIbh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2rxIbh_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.stateTable2rxIbh_rsp_U' read by process 'rocev2_top_rocev2_top.state_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.stateTable2rxIbh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    22: begin
                        if (~rx_ibh_fsm_0_U0.rx_ibhDropFifo_blk_n) begin
                            if (~rx_ibhDropFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibhDropFifo_U' written by process 'rocev2_top_rocev2_top.drop_ooo_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhDropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibhDropFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibhDropFifo_U' read by process 'rocev2_top_rocev2_top.drop_ooo_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhDropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    23: begin
                        if (~rx_ibh_fsm_0_U0.rx_ibhDropMetaFifo_blk_n) begin
                            if (~rx_ibhDropMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibhDropMetaFifo_U' written by process 'rocev2_top_rocev2_top.ipUdpMetaHandler_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhDropMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibhDropMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibhDropMetaFifo_U' read by process 'rocev2_top_rocev2_top.ipUdpMetaHandler_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhDropMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    24: begin
                        if (~rx_ibh_fsm_0_U0.rx_fsm2exh_MetaFifo_blk_n) begin
                            if (~rx_fsm2exh_MetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_fsm2exh_MetaFifo_U' written by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_fsm2exh_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_fsm2exh_MetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_fsm2exh_MetaFifo_U' read by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_fsm2exh_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    51: begin
                        if (~rx_ibh_fsm_0_U0.rx2retrans_upd_blk_n) begin
                            if (~rx2retrans_upd_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx2retrans_upd_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx2retrans_upd_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx2retrans_upd_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx2retrans_upd_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx2retrans_upd_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    47: begin
                        if (~rx_ibh_fsm_0_U0.rxClearTimer_req_blk_n) begin
                            if (~rxClearTimer_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rxClearTimer_req_U' written by process 'rocev2_top_rocev2_top.transport_timer_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rxClearTimer_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxClearTimer_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rxClearTimer_req_U' read by process 'rocev2_top_rocev2_top.transport_timer_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rxClearTimer_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    27: begin
                        if (~rx_ibh_fsm_0_U0.rx_ibhEventFifo_blk_n) begin
                            if (~rx_ibhEventFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibhEventFifo_U' written by process 'rocev2_top_rocev2_top.stream_merger_ackEvent_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibhEventFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibhEventFifo_U' read by process 'rocev2_top_rocev2_top.stream_merger_ackEvent_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                22 : begin
                    case(index2)
                    21: begin
                        if (~drop_ooo_ibh_512_0_U0.rx_ibhDropFifo_blk_n) begin
                            if (~rx_ibhDropFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibhDropFifo_U' written by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhDropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibhDropFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibhDropFifo_U' read by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhDropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (~drop_ooo_ibh_512_0_U0.rx_exh2dropFifo_blk_n) begin
                            if (~rx_exh2dropFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exh2dropFifo_U' written by process 'rocev2_top_rocev2_top.rx_process_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2dropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exh2dropFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exh2dropFifo_U' read by process 'rocev2_top_rocev2_top.rx_process_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2dropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    25: begin
                        if (~drop_ooo_ibh_512_0_U0.rx_ibhDrop2exhFifo_blk_n) begin
                            if (~rx_ibhDrop2exhFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibhDrop2exhFifo_U' written by process 'rocev2_top_rocev2_top.rx_exh_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhDrop2exhFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibhDrop2exhFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibhDrop2exhFifo_U' read by process 'rocev2_top_rocev2_top.rx_exh_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhDrop2exhFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                23 : begin
                    case(index2)
                    13: begin
                        if (~ipUdpMetaHandler_512_0_U0.rx_ipUdpMetaFifo_blk_n) begin
                            if (~rx_ipUdpMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ipUdpMetaFifo_U' written by process 'rocev2_top_rocev2_top.merge_rx_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ipUdpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ipUdpMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ipUdpMetaFifo_U' read by process 'rocev2_top_rocev2_top.merge_rx_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ipUdpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (~ipUdpMetaHandler_512_0_U0.rx_exh2drop_MetaFifo_blk_n) begin
                            if (~rx_exh2drop_MetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exh2drop_MetaFifo_U' written by process 'rocev2_top_rocev2_top.rx_process_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2drop_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exh2drop_MetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exh2drop_MetaFifo_U' read by process 'rocev2_top_rocev2_top.rx_process_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2drop_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    21: begin
                        if (~ipUdpMetaHandler_512_0_U0.rx_ibhDropMetaFifo_blk_n) begin
                            if (~rx_ibhDropMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibhDropMetaFifo_U' written by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhDropMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibhDropMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibhDropMetaFifo_U' read by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhDropMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    24: begin
                        if (~ipUdpMetaHandler_512_0_U0.exh_lengthFifo_blk_n) begin
                            if (~exh_lengthFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.exh_lengthFifo_U' written by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.exh_lengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~exh_lengthFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.exh_lengthFifo_U' read by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.exh_lengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~ipUdpMetaHandler_512_0_U0.rx_drop2exhFsm_MetaFifo_blk_n) begin
                            if (~rx_drop2exhFsm_MetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_drop2exhFsm_MetaFifo_U' written by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_drop2exhFsm_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_drop2exhFsm_MetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_drop2exhFsm_MetaFifo_U' read by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_drop2exhFsm_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                24 : begin
                    case(index2)
                    21: begin
                        if (~rx_exh_fsm_512_0_U0.rx_fsm2exh_MetaFifo_blk_n) begin
                            if (~rx_fsm2exh_MetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_fsm2exh_MetaFifo_U' written by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_fsm2exh_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_fsm2exh_MetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_fsm2exh_MetaFifo_U' read by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_fsm2exh_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    23: begin
                        if (~rx_exh_fsm_512_0_U0.rx_drop2exhFsm_MetaFifo_blk_n) begin
                            if (~rx_drop2exhFsm_MetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_drop2exhFsm_MetaFifo_U' written by process 'rocev2_top_rocev2_top.ipUdpMetaHandler_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_drop2exhFsm_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_drop2exhFsm_MetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_drop2exhFsm_MetaFifo_U' read by process 'rocev2_top_rocev2_top.ipUdpMetaHandler_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_drop2exhFsm_MetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rx_exh_fsm_512_0_U0.exh_lengthFifo_blk_n) begin
                            if (~exh_lengthFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.exh_lengthFifo_U' written by process 'rocev2_top_rocev2_top.ipUdpMetaHandler_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.exh_lengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~exh_lengthFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.exh_lengthFifo_U' read by process 'rocev2_top_rocev2_top.ipUdpMetaHandler_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.exh_lengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    45: begin
                        if (~rx_exh_fsm_512_0_U0.rxExh2msnTable_upd_req_blk_n) begin
                            if (~rxExh2msnTable_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rxExh2msnTable_upd_req_U' written by process 'rocev2_top_rocev2_top.msn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rxExh2msnTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxExh2msnTable_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rxExh2msnTable_upd_req_U' read by process 'rocev2_top_rocev2_top.msn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rxExh2msnTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rx_exh_fsm_512_0_U0.msnTable2rxExh_rsp_blk_n) begin
                            if (~msnTable2rxExh_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.msnTable2rxExh_rsp_U' written by process 'rocev2_top_rocev2_top.msn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.msnTable2rxExh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~msnTable2rxExh_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.msnTable2rxExh_rsp_U' read by process 'rocev2_top_rocev2_top.msn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.msnTable2rxExh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    51: begin
                        if (~rx_exh_fsm_512_0_U0.retrans2rx_init_blk_n) begin
                            if (~retrans2rx_init_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.retrans2rx_init_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.retrans2rx_init_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~retrans2rx_init_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.retrans2rx_init_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.retrans2rx_init_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rx_exh_fsm_512_0_U0.rx2retrans_req_blk_n) begin
                            if (~rx2retrans_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx2retrans_req_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx2retrans_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx2retrans_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx2retrans_req_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx2retrans_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    27: begin
                        if (~rx_exh_fsm_512_0_U0.rx_exhEventMetaFifo_blk_n) begin
                            if (~rx_exhEventMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exhEventMetaFifo_U' written by process 'rocev2_top_rocev2_top.stream_merger_ackEvent_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exhEventMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exhEventMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exhEventMetaFifo_U' read by process 'rocev2_top_rocev2_top.stream_merger_ackEvent_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exhEventMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    25: begin
                        if (~rx_exh_fsm_512_0_U0.rx_pkgSplitTypeFifo_blk_n) begin
                            if (~rx_pkgSplitTypeFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_pkgSplitTypeFifo_U' written by process 'rocev2_top_rocev2_top.rx_exh_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_pkgSplitTypeFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_pkgSplitTypeFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_pkgSplitTypeFifo_U' read by process 'rocev2_top_rocev2_top.rx_exh_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_pkgSplitTypeFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    30: begin
                        if (~rx_exh_fsm_512_0_U0.rx_pkgShiftTypeFifo_blk_n) begin
                            if (~rx_pkgShiftTypeFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_pkgShiftTypeFifo_U' written by process 'rocev2_top_rocev2_top.merge_rx_pkgs_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_pkgShiftTypeFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_pkgShiftTypeFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_pkgShiftTypeFifo_U' read by process 'rocev2_top_rocev2_top.merge_rx_pkgs_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_pkgShiftTypeFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    26: begin
                        if (~rx_exh_fsm_512_0_U0.rx_readRequestFifo_blk_n) begin
                            if (~rx_readRequestFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_readRequestFifo_U' written by process 'rocev2_top_rocev2_top.handle_read_requests_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_readRequestFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_readRequestFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_readRequestFifo_U' read by process 'rocev2_top_rocev2_top.handle_read_requests_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_readRequestFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                25 : begin
                    case(index2)
                    24: begin
                        if (~rx_exh_payload_512_0_U0.rx_pkgSplitTypeFifo_blk_n) begin
                            if (~rx_pkgSplitTypeFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_pkgSplitTypeFifo_U' written by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_pkgSplitTypeFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_pkgSplitTypeFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_pkgSplitTypeFifo_U' read by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_pkgSplitTypeFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    22: begin
                        if (~rx_exh_payload_512_0_U0.rx_ibhDrop2exhFifo_blk_n) begin
                            if (~rx_ibhDrop2exhFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibhDrop2exhFifo_U' written by process 'rocev2_top_rocev2_top.drop_ooo_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhDrop2exhFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibhDrop2exhFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibhDrop2exhFifo_U' read by process 'rocev2_top_rocev2_top.drop_ooo_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhDrop2exhFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    28: begin
                        if (~rx_exh_payload_512_0_U0.rx_exh2rethShiftFifo_blk_n) begin
                            if (~rx_exh2rethShiftFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exh2rethShiftFifo_U' written by process 'rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_12_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2rethShiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exh2rethShiftFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exh2rethShiftFifo_U' read by process 'rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_12_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2rethShiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    29: begin
                        if (~rx_exh_payload_512_0_U0.rx_exh2aethShiftFifo_blk_n) begin
                            if (~rx_exh2aethShiftFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exh2aethShiftFifo_U' written by process 'rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_13_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2aethShiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exh2aethShiftFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exh2aethShiftFifo_U' read by process 'rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_13_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2aethShiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    30: begin
                        if (~rx_exh_payload_512_0_U0.rx_exhNoShiftFifo_blk_n) begin
                            if (~rx_exhNoShiftFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exhNoShiftFifo_U' written by process 'rocev2_top_rocev2_top.merge_rx_pkgs_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exhNoShiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exhNoShiftFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exhNoShiftFifo_U' read by process 'rocev2_top_rocev2_top.merge_rx_pkgs_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exhNoShiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                26 : begin
                    case(index2)
                    24: begin
                        if (~handle_read_requests_0_U0.rx_readRequestFifo_blk_n) begin
                            if (~rx_readRequestFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_readRequestFifo_U' written by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_readRequestFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_readRequestFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_readRequestFifo_U' read by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_readRequestFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    42: begin
                        if (~handle_read_requests_0_U0.rx_remoteMemCmd_blk_n) begin
                            if (~rx_remoteMemCmd_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_remoteMemCmd_U' written by process 'rocev2_top_rocev2_top.mem_cmd_merger_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_remoteMemCmd_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_remoteMemCmd_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_remoteMemCmd_U' read by process 'rocev2_top_rocev2_top.mem_cmd_merger_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_remoteMemCmd_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    33: begin
                        if (~handle_read_requests_0_U0.rx_readEvenFifo_blk_n) begin
                            if (~rx_readEvenFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_readEvenFifo_U' written by process 'rocev2_top_rocev2_top.meta_merger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_readEvenFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_readEvenFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_readEvenFifo_U' read by process 'rocev2_top_rocev2_top.meta_merger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_readEvenFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                27 : begin
                    case(index2)
                    24: begin
                        if (~stream_merger_ackEvent_U0.rx_exhEventMetaFifo_blk_n) begin
                            if (~rx_exhEventMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exhEventMetaFifo_U' written by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exhEventMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exhEventMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exhEventMetaFifo_U' read by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exhEventMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    33: begin
                        if (~stream_merger_ackEvent_U0.rx_ackEventFifo_blk_n) begin
                            if (~rx_ackEventFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ackEventFifo_U' written by process 'rocev2_top_rocev2_top.meta_merger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ackEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ackEventFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ackEventFifo_U' read by process 'rocev2_top_rocev2_top.meta_merger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ackEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    21: begin
                        if (~stream_merger_ackEvent_U0.rx_ibhEventFifo_blk_n) begin
                            if (~rx_ibhEventFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ibhEventFifo_U' written by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ibhEventFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ibhEventFifo_U' read by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ibhEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                28 : begin
                    case(index2)
                    25: begin
                        if (~rshiftWordByOctet_net_axis_512_512_12_0_U0.rx_exh2rethShiftFifo_blk_n) begin
                            if (~rx_exh2rethShiftFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exh2rethShiftFifo_U' written by process 'rocev2_top_rocev2_top.rx_exh_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2rethShiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exh2rethShiftFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exh2rethShiftFifo_U' read by process 'rocev2_top_rocev2_top.rx_exh_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2rethShiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    30: begin
                        if (~rshiftWordByOctet_net_axis_512_512_12_0_U0.rx_rethSift2mergerFifo_blk_n) begin
                            if (~rx_rethSift2mergerFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_rethSift2mergerFifo_U' written by process 'rocev2_top_rocev2_top.merge_rx_pkgs_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_rethSift2mergerFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_rethSift2mergerFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_rethSift2mergerFifo_U' read by process 'rocev2_top_rocev2_top.merge_rx_pkgs_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_rethSift2mergerFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                29 : begin
                    case(index2)
                    25: begin
                        if (~rshiftWordByOctet_net_axis_512_512_13_0_U0.rx_exh2aethShiftFifo_blk_n) begin
                            if (~rx_exh2aethShiftFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exh2aethShiftFifo_U' written by process 'rocev2_top_rocev2_top.rx_exh_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2aethShiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exh2aethShiftFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exh2aethShiftFifo_U' read by process 'rocev2_top_rocev2_top.rx_exh_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exh2aethShiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    30: begin
                        if (~rshiftWordByOctet_net_axis_512_512_13_0_U0.rx_aethSift2mergerFifo_blk_n) begin
                            if (~rx_aethSift2mergerFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_aethSift2mergerFifo_U' written by process 'rocev2_top_rocev2_top.merge_rx_pkgs_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_aethSift2mergerFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_aethSift2mergerFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_aethSift2mergerFifo_U' read by process 'rocev2_top_rocev2_top.merge_rx_pkgs_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_aethSift2mergerFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                30 : begin
                    case(index2)
                    24: begin
                        if (~merge_rx_pkgs_512_0_U0.rx_pkgShiftTypeFifo_blk_n) begin
                            if (~rx_pkgShiftTypeFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_pkgShiftTypeFifo_U' written by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_pkgShiftTypeFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_pkgShiftTypeFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_pkgShiftTypeFifo_U' read by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_pkgShiftTypeFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    29: begin
                        if (~merge_rx_pkgs_512_0_U0.rx_aethSift2mergerFifo_blk_n) begin
                            if (~rx_aethSift2mergerFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_aethSift2mergerFifo_U' written by process 'rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_13_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_aethSift2mergerFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_aethSift2mergerFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_aethSift2mergerFifo_U' read by process 'rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_13_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_aethSift2mergerFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    4: begin
                        if (~merge_rx_pkgs_512_0_U0.m_axis_mem_write_data_internal_blk_n) begin
                            if (~m_axis_mem_write_data_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.m_axis_mem_write_data_internal_U' written by process 'rocev2_top_rocev2_top.convert_net_axis_to_axis_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.m_axis_mem_write_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~m_axis_mem_write_data_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.m_axis_mem_write_data_internal_U' read by process 'rocev2_top_rocev2_top.convert_net_axis_to_axis_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.m_axis_mem_write_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    28: begin
                        if (~merge_rx_pkgs_512_0_U0.rx_rethSift2mergerFifo_blk_n) begin
                            if (~rx_rethSift2mergerFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_rethSift2mergerFifo_U' written by process 'rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_12_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_rethSift2mergerFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_rethSift2mergerFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_rethSift2mergerFifo_U' read by process 'rocev2_top_rocev2_top.rshiftWordByOctet_net_axis_512_512_12_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_rethSift2mergerFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    25: begin
                        if (~merge_rx_pkgs_512_0_U0.rx_exhNoShiftFifo_blk_n) begin
                            if (~rx_exhNoShiftFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_exhNoShiftFifo_U' written by process 'rocev2_top_rocev2_top.rx_exh_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exhNoShiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_exhNoShiftFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_exhNoShiftFifo_U' read by process 'rocev2_top_rocev2_top.rx_exh_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_exhNoShiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                31 : begin
                    case(index2)
                    51: begin
                        if (~local_req_handler_0_U0.retransmitter2exh_eventFifo_blk_n) begin
                            if (~retransmitter2exh_eventFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.retransmitter2exh_eventFifo_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.retransmitter2exh_eventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~retransmitter2exh_eventFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.retransmitter2exh_eventFifo_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.retransmitter2exh_eventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    33: begin
                        if (~local_req_handler_0_U0.tx_appMetaFifo_blk_n) begin
                            if (~tx_appMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_appMetaFifo_U' written by process 'rocev2_top_rocev2_top.meta_merger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_appMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_appMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_appMetaFifo_U' read by process 'rocev2_top_rocev2_top.meta_merger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_appMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    42: begin
                        if (~local_req_handler_0_U0.tx_localMemCmdFifo_blk_n) begin
                            if (~tx_localMemCmdFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_localMemCmdFifo_U' written by process 'rocev2_top_rocev2_top.mem_cmd_merger_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_localMemCmdFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_localMemCmdFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_localMemCmdFifo_U' read by process 'rocev2_top_rocev2_top.mem_cmd_merger_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_localMemCmdFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    46: begin
                        if (~local_req_handler_0_U0.tx2retrans_insertAddrLen_blk_n) begin
                            if (~tx2retrans_insertAddrLen_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx2retrans_insertAddrLen_U' written by process 'rocev2_top_rocev2_top.merge_retrans_request_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx2retrans_insertAddrLen_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx2retrans_insertAddrLen_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx2retrans_insertAddrLen_U' read by process 'rocev2_top_rocev2_top.merge_retrans_request_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx2retrans_insertAddrLen_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                32 : begin
                    case(index2)
                    42: begin
                        if (~tx_pkg_arbiter_512_0_U0.tx_pkgInfoFifo_blk_n) begin
                            if (~tx_pkgInfoFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_pkgInfoFifo_U' written by process 'rocev2_top_rocev2_top.mem_cmd_merger_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_pkgInfoFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_pkgInfoFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_pkgInfoFifo_U' read by process 'rocev2_top_rocev2_top.mem_cmd_merger_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_pkgInfoFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    3: begin
                        if (~tx_pkg_arbiter_512_0_U0.s_axis_mem_read_data_internal_blk_n) begin
                            if (~s_axis_mem_read_data_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.s_axis_mem_read_data_internal_U' written by process 'rocev2_top_rocev2_top.convert_axis_to_net_axis_512_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.s_axis_mem_read_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~s_axis_mem_read_data_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.s_axis_mem_read_data_internal_U' read by process 'rocev2_top_rocev2_top.convert_axis_to_net_axis_512_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.s_axis_mem_read_data_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    34: begin
                        if (~tx_pkg_arbiter_512_0_U0.tx_split2aethShift_blk_n) begin
                            if (~tx_split2aethShift_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_split2aethShift_U' written by process 'rocev2_top_rocev2_top.lshiftWordByOctet_512_12_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_split2aethShift_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_split2aethShift_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_split2aethShift_U' read by process 'rocev2_top_rocev2_top.lshiftWordByOctet_512_12_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_split2aethShift_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    35: begin
                        if (~tx_pkg_arbiter_512_0_U0.tx_rethMerge2rethShift_blk_n) begin
                            if (~tx_rethMerge2rethShift_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_rethMerge2rethShift_U' written by process 'rocev2_top_rocev2_top.lshiftWordByOctet_512_13_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_rethMerge2rethShift_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_rethMerge2rethShift_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_rethMerge2rethShift_U' read by process 'rocev2_top_rocev2_top.lshiftWordByOctet_512_13_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_rethMerge2rethShift_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    37: begin
                        if (~tx_pkg_arbiter_512_0_U0.tx_rawPayFifo_blk_n) begin
                            if (~tx_rawPayFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_rawPayFifo_U' written by process 'rocev2_top_rocev2_top.append_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_rawPayFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_rawPayFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_rawPayFifo_U' read by process 'rocev2_top_rocev2_top.append_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_rawPayFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                33 : begin
                    case(index2)
                    27: begin
                        if (~meta_merger_0_U0.rx_ackEventFifo_blk_n) begin
                            if (~rx_ackEventFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_ackEventFifo_U' written by process 'rocev2_top_rocev2_top.stream_merger_ackEvent_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ackEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_ackEventFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_ackEventFifo_U' read by process 'rocev2_top_rocev2_top.stream_merger_ackEvent_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_ackEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    43: begin
                        if (~meta_merger_0_U0.tx_ibhconnTable_req_blk_n) begin
                            if (~tx_ibhconnTable_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_ibhconnTable_req_U' written by process 'rocev2_top_rocev2_top.conn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ibhconnTable_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_ibhconnTable_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_ibhconnTable_req_U' read by process 'rocev2_top_rocev2_top.conn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ibhconnTable_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    39: begin
                        if (~meta_merger_0_U0.tx_ibhMetaFifo_blk_n) begin
                            if (~tx_ibhMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_ibhMetaFifo_U' written by process 'rocev2_top_rocev2_top.generate_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ibhMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_ibhMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_ibhMetaFifo_U' read by process 'rocev2_top_rocev2_top.generate_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ibhMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    36: begin
                        if (~meta_merger_0_U0.tx_exhMetaFifo_blk_n) begin
                            if (~tx_exhMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_exhMetaFifo_U' written by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_exhMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_exhMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_exhMetaFifo_U' read by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_exhMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    26: begin
                        if (~meta_merger_0_U0.rx_readEvenFifo_blk_n) begin
                            if (~rx_readEvenFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_readEvenFifo_U' written by process 'rocev2_top_rocev2_top.handle_read_requests_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_readEvenFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_readEvenFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_readEvenFifo_U' read by process 'rocev2_top_rocev2_top.handle_read_requests_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_readEvenFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    31: begin
                        if (~meta_merger_0_U0.tx_appMetaFifo_blk_n) begin
                            if (~tx_appMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_appMetaFifo_U' written by process 'rocev2_top_rocev2_top.local_req_handler_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_appMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_appMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_appMetaFifo_U' read by process 'rocev2_top_rocev2_top.local_req_handler_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_appMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                34 : begin
                    case(index2)
                    37: begin
                        if (~lshiftWordByOctet_512_12_0_U0.tx_aethShift2payFifo_blk_n) begin
                            if (~tx_aethShift2payFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_aethShift2payFifo_U' written by process 'rocev2_top_rocev2_top.append_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_aethShift2payFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_aethShift2payFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_aethShift2payFifo_U' read by process 'rocev2_top_rocev2_top.append_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_aethShift2payFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    32: begin
                        if (~lshiftWordByOctet_512_12_0_U0.tx_split2aethShift_blk_n) begin
                            if (~tx_split2aethShift_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_split2aethShift_U' written by process 'rocev2_top_rocev2_top.tx_pkg_arbiter_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_split2aethShift_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_split2aethShift_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_split2aethShift_U' read by process 'rocev2_top_rocev2_top.tx_pkg_arbiter_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_split2aethShift_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                35 : begin
                    case(index2)
                    37: begin
                        if (~lshiftWordByOctet_512_13_0_U0.tx_rethShift2payFifo_blk_n) begin
                            if (~tx_rethShift2payFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_rethShift2payFifo_U' written by process 'rocev2_top_rocev2_top.append_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_rethShift2payFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_rethShift2payFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_rethShift2payFifo_U' read by process 'rocev2_top_rocev2_top.append_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_rethShift2payFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    32: begin
                        if (~lshiftWordByOctet_512_13_0_U0.tx_rethMerge2rethShift_blk_n) begin
                            if (~tx_rethMerge2rethShift_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_rethMerge2rethShift_U' written by process 'rocev2_top_rocev2_top.tx_pkg_arbiter_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_rethMerge2rethShift_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_rethMerge2rethShift_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_rethMerge2rethShift_U' read by process 'rocev2_top_rocev2_top.tx_pkg_arbiter_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_rethMerge2rethShift_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                36 : begin
                    case(index2)
                    33: begin
                        if (~generate_exh_512_0_U0.tx_exhMetaFifo_blk_n) begin
                            if (~tx_exhMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_exhMetaFifo_U' written by process 'rocev2_top_rocev2_top.meta_merger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_exhMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_exhMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_exhMetaFifo_U' read by process 'rocev2_top_rocev2_top.meta_merger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_exhMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    45: begin
                        if (~generate_exh_512_0_U0.txExh2msnTable_req_blk_n) begin
                            if (~txExh2msnTable_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.txExh2msnTable_req_U' written by process 'rocev2_top_rocev2_top.msn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.txExh2msnTable_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txExh2msnTable_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.txExh2msnTable_req_U' read by process 'rocev2_top_rocev2_top.msn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.txExh2msnTable_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~generate_exh_512_0_U0.msnTable2txExh_rsp_blk_n) begin
                            if (~msnTable2txExh_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.msnTable2txExh_rsp_U' written by process 'rocev2_top_rocev2_top.msn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.msnTable2txExh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~msnTable2txExh_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.msnTable2txExh_rsp_U' read by process 'rocev2_top_rocev2_top.msn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.msnTable2txExh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    47: begin
                        if (~generate_exh_512_0_U0.txSetTimer_req_blk_n) begin
                            if (~txSetTimer_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.txSetTimer_req_U' written by process 'rocev2_top_rocev2_top.transport_timer_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.txSetTimer_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txSetTimer_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.txSetTimer_req_U' read by process 'rocev2_top_rocev2_top.transport_timer_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.txSetTimer_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    37: begin
                        if (~generate_exh_512_0_U0.tx_exh2payFifo_blk_n) begin
                            if (~tx_exh2payFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_exh2payFifo_U' written by process 'rocev2_top_rocev2_top.append_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_exh2payFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_exh2payFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_exh2payFifo_U' read by process 'rocev2_top_rocev2_top.append_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_exh2payFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~generate_exh_512_0_U0.tx_packetInfoFifo_blk_n) begin
                            if (~tx_packetInfoFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_packetInfoFifo_U' written by process 'rocev2_top_rocev2_top.append_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_packetInfoFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_packetInfoFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_packetInfoFifo_U' read by process 'rocev2_top_rocev2_top.append_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_packetInfoFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    41: begin
                        if (~generate_exh_512_0_U0.tx_lengthFifo_blk_n) begin
                            if (~tx_lengthFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_lengthFifo_U' written by process 'rocev2_top_rocev2_top.tx_ipUdpMetaMerger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_lengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_lengthFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_lengthFifo_U' read by process 'rocev2_top_rocev2_top.tx_ipUdpMetaMerger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_lengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                37 : begin
                    case(index2)
                    36: begin
                        if (~append_payload_512_0_U0.tx_packetInfoFifo_blk_n) begin
                            if (~tx_packetInfoFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_packetInfoFifo_U' written by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_packetInfoFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_packetInfoFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_packetInfoFifo_U' read by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_packetInfoFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~append_payload_512_0_U0.tx_exh2payFifo_blk_n) begin
                            if (~tx_exh2payFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_exh2payFifo_U' written by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_exh2payFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_exh2payFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_exh2payFifo_U' read by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_exh2payFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    38: begin
                        if (~append_payload_512_0_U0.tx_exh2shiftFifo_blk_n) begin
                            if (~tx_exh2shiftFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_exh2shiftFifo_U' written by process 'rocev2_top_rocev2_top.lshiftWordByOctet_512_11_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_exh2shiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_exh2shiftFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_exh2shiftFifo_U' read by process 'rocev2_top_rocev2_top.lshiftWordByOctet_512_11_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_exh2shiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    34: begin
                        if (~append_payload_512_0_U0.tx_aethShift2payFifo_blk_n) begin
                            if (~tx_aethShift2payFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_aethShift2payFifo_U' written by process 'rocev2_top_rocev2_top.lshiftWordByOctet_512_12_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_aethShift2payFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_aethShift2payFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_aethShift2payFifo_U' read by process 'rocev2_top_rocev2_top.lshiftWordByOctet_512_12_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_aethShift2payFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    35: begin
                        if (~append_payload_512_0_U0.tx_rethShift2payFifo_blk_n) begin
                            if (~tx_rethShift2payFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_rethShift2payFifo_U' written by process 'rocev2_top_rocev2_top.lshiftWordByOctet_512_13_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_rethShift2payFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_rethShift2payFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_rethShift2payFifo_U' read by process 'rocev2_top_rocev2_top.lshiftWordByOctet_512_13_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_rethShift2payFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    32: begin
                        if (~append_payload_512_0_U0.tx_rawPayFifo_blk_n) begin
                            if (~tx_rawPayFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_rawPayFifo_U' written by process 'rocev2_top_rocev2_top.tx_pkg_arbiter_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_rawPayFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_rawPayFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_rawPayFifo_U' read by process 'rocev2_top_rocev2_top.tx_pkg_arbiter_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_rawPayFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                38 : begin
                    case(index2)
                    40: begin
                        if (~lshiftWordByOctet_512_11_0_U0.tx_shift2ibhFifo_blk_n) begin
                            if (~tx_shift2ibhFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_shift2ibhFifo_U' written by process 'rocev2_top_rocev2_top.prepend_ibh_header_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_shift2ibhFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_shift2ibhFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_shift2ibhFifo_U' read by process 'rocev2_top_rocev2_top.prepend_ibh_header_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_shift2ibhFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    37: begin
                        if (~lshiftWordByOctet_512_11_0_U0.tx_exh2shiftFifo_blk_n) begin
                            if (~tx_exh2shiftFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_exh2shiftFifo_U' written by process 'rocev2_top_rocev2_top.append_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_exh2shiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_exh2shiftFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_exh2shiftFifo_U' read by process 'rocev2_top_rocev2_top.append_payload_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_exh2shiftFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                39 : begin
                    case(index2)
                    33: begin
                        if (~generate_ibh_512_0_U0.tx_ibhMetaFifo_blk_n) begin
                            if (~tx_ibhMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_ibhMetaFifo_U' written by process 'rocev2_top_rocev2_top.meta_merger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ibhMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_ibhMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_ibhMetaFifo_U' read by process 'rocev2_top_rocev2_top.meta_merger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ibhMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    41: begin
                        if (~generate_ibh_512_0_U0.tx_dstQpFifo_blk_n) begin
                            if (~tx_dstQpFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_dstQpFifo_U' written by process 'rocev2_top_rocev2_top.tx_ipUdpMetaMerger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_dstQpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_dstQpFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_dstQpFifo_U' read by process 'rocev2_top_rocev2_top.tx_ipUdpMetaMerger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_dstQpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    40: begin
                        if (~generate_ibh_512_0_U0.tx_ibhHeaderFifo_blk_n) begin
                            if (~tx_ibhHeaderFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_ibhHeaderFifo_U' written by process 'rocev2_top_rocev2_top.prepend_ibh_header_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ibhHeaderFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_ibhHeaderFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_ibhHeaderFifo_U' read by process 'rocev2_top_rocev2_top.prepend_ibh_header_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ibhHeaderFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    44: begin
                        if (~generate_ibh_512_0_U0.txIbh2stateTable_upd_req_blk_n) begin
                            if (~txIbh2stateTable_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.txIbh2stateTable_upd_req_U' written by process 'rocev2_top_rocev2_top.state_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.txIbh2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txIbh2stateTable_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.txIbh2stateTable_upd_req_U' read by process 'rocev2_top_rocev2_top.state_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.txIbh2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~generate_ibh_512_0_U0.stateTable2txIbh_rsp_blk_n) begin
                            if (~stateTable2txIbh_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.stateTable2txIbh_rsp_U' written by process 'rocev2_top_rocev2_top.state_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.stateTable2txIbh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2txIbh_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.stateTable2txIbh_rsp_U' read by process 'rocev2_top_rocev2_top.state_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.stateTable2txIbh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    46: begin
                        if (~generate_ibh_512_0_U0.tx2retrans_insertMeta_blk_n) begin
                            if (~tx2retrans_insertMeta_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx2retrans_insertMeta_U' written by process 'rocev2_top_rocev2_top.merge_retrans_request_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx2retrans_insertMeta_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx2retrans_insertMeta_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx2retrans_insertMeta_U' read by process 'rocev2_top_rocev2_top.merge_retrans_request_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx2retrans_insertMeta_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                40 : begin
                    case(index2)
                    39: begin
                        if (~prepend_ibh_header_512_0_U0.tx_ibhHeaderFifo_blk_n) begin
                            if (~tx_ibhHeaderFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_ibhHeaderFifo_U' written by process 'rocev2_top_rocev2_top.generate_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ibhHeaderFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_ibhHeaderFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_ibhHeaderFifo_U' read by process 'rocev2_top_rocev2_top.generate_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ibhHeaderFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    15: begin
                        if (~prepend_ibh_header_512_0_U0.tx_ib2udpFifo_blk_n) begin
                            if (~tx_ib2udpFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_ib2udpFifo_U' written by process 'rocev2_top_rocev2_top.udp_lshiftWordByOctet_512_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ib2udpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_ib2udpFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_ib2udpFifo_U' read by process 'rocev2_top_rocev2_top.udp_lshiftWordByOctet_512_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ib2udpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    38: begin
                        if (~prepend_ibh_header_512_0_U0.tx_shift2ibhFifo_blk_n) begin
                            if (~tx_shift2ibhFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_shift2ibhFifo_U' written by process 'rocev2_top_rocev2_top.lshiftWordByOctet_512_11_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_shift2ibhFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_shift2ibhFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_shift2ibhFifo_U' read by process 'rocev2_top_rocev2_top.lshiftWordByOctet_512_11_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_shift2ibhFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                41 : begin
                    case(index2)
                    43: begin
                        if (~tx_ipUdpMetaMerger_0_U0.tx_connTable2ibh_rsp_blk_n) begin
                            if (~tx_connTable2ibh_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_connTable2ibh_rsp_U' written by process 'rocev2_top_rocev2_top.conn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_connTable2ibh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_connTable2ibh_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_connTable2ibh_rsp_U' read by process 'rocev2_top_rocev2_top.conn_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_connTable2ibh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    36: begin
                        if (~tx_ipUdpMetaMerger_0_U0.tx_lengthFifo_blk_n) begin
                            if (~tx_lengthFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_lengthFifo_U' written by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_lengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_lengthFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_lengthFifo_U' read by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_lengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (~tx_ipUdpMetaMerger_0_U0.tx_ipUdpMetaFifo_blk_n) begin
                            if (~tx_ipUdpMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_ipUdpMetaFifo_U' written by process 'rocev2_top_rocev2_top.split_tx_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ipUdpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_ipUdpMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_ipUdpMetaFifo_U' read by process 'rocev2_top_rocev2_top.split_tx_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ipUdpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    39: begin
                        if (~tx_ipUdpMetaMerger_0_U0.tx_dstQpFifo_blk_n) begin
                            if (~tx_dstQpFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_dstQpFifo_U' written by process 'rocev2_top_rocev2_top.generate_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_dstQpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_dstQpFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_dstQpFifo_U' read by process 'rocev2_top_rocev2_top.generate_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_dstQpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                42 : begin
                    case(index2)
                    26: begin
                        if (~mem_cmd_merger_512_0_U0.rx_remoteMemCmd_blk_n) begin
                            if (~rx_remoteMemCmd_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx_remoteMemCmd_U' written by process 'rocev2_top_rocev2_top.handle_read_requests_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_remoteMemCmd_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_remoteMemCmd_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx_remoteMemCmd_U' read by process 'rocev2_top_rocev2_top.handle_read_requests_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx_remoteMemCmd_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    32: begin
                        if (~mem_cmd_merger_512_0_U0.tx_pkgInfoFifo_blk_n) begin
                            if (~tx_pkgInfoFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_pkgInfoFifo_U' written by process 'rocev2_top_rocev2_top.tx_pkg_arbiter_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_pkgInfoFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_pkgInfoFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_pkgInfoFifo_U' read by process 'rocev2_top_rocev2_top.tx_pkg_arbiter_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_pkgInfoFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    31: begin
                        if (~mem_cmd_merger_512_0_U0.tx_localMemCmdFifo_blk_n) begin
                            if (~tx_localMemCmdFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_localMemCmdFifo_U' written by process 'rocev2_top_rocev2_top.local_req_handler_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_localMemCmdFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_localMemCmdFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_localMemCmdFifo_U' read by process 'rocev2_top_rocev2_top.local_req_handler_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_localMemCmdFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                43 : begin
                    case(index2)
                    33: begin
                        if (~conn_table_0_U0.tx_ibhconnTable_req_blk_n) begin
                            if (~tx_ibhconnTable_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_ibhconnTable_req_U' written by process 'rocev2_top_rocev2_top.meta_merger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ibhconnTable_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_ibhconnTable_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_ibhconnTable_req_U' read by process 'rocev2_top_rocev2_top.meta_merger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_ibhconnTable_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    41: begin
                        if (~conn_table_0_U0.tx_connTable2ibh_rsp_blk_n) begin
                            if (~tx_connTable2ibh_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx_connTable2ibh_rsp_U' written by process 'rocev2_top_rocev2_top.tx_ipUdpMetaMerger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_connTable2ibh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx_connTable2ibh_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx_connTable2ibh_rsp_U' read by process 'rocev2_top_rocev2_top.tx_ipUdpMetaMerger_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx_connTable2ibh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                44 : begin
                    case(index2)
                    21: begin
                        if (~state_table_0_U0.rxIbh2stateTable_upd_req_blk_n) begin
                            if (~rxIbh2stateTable_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rxIbh2stateTable_upd_req_U' written by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rxIbh2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxIbh2stateTable_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rxIbh2stateTable_upd_req_U' read by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rxIbh2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~state_table_0_U0.stateTable2rxIbh_rsp_blk_n) begin
                            if (~stateTable2rxIbh_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.stateTable2rxIbh_rsp_U' written by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.stateTable2rxIbh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2rxIbh_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.stateTable2rxIbh_rsp_U' read by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.stateTable2rxIbh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    39: begin
                        if (~state_table_0_U0.txIbh2stateTable_upd_req_blk_n) begin
                            if (~txIbh2stateTable_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.txIbh2stateTable_upd_req_U' written by process 'rocev2_top_rocev2_top.generate_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.txIbh2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txIbh2stateTable_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.txIbh2stateTable_upd_req_U' read by process 'rocev2_top_rocev2_top.generate_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.txIbh2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~state_table_0_U0.stateTable2txIbh_rsp_blk_n) begin
                            if (~stateTable2txIbh_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.stateTable2txIbh_rsp_U' written by process 'rocev2_top_rocev2_top.generate_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.stateTable2txIbh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2txIbh_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.stateTable2txIbh_rsp_U' read by process 'rocev2_top_rocev2_top.generate_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.stateTable2txIbh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    17: begin
                        if (~state_table_0_U0.qpi2stateTable_upd_req_blk_n) begin
                            if (~qpi2stateTable_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.qpi2stateTable_upd_req_U' written by process 'rocev2_top_rocev2_top.qp_interface_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.qpi2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~qpi2stateTable_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.qpi2stateTable_upd_req_U' read by process 'rocev2_top_rocev2_top.qp_interface_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.qpi2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~state_table_0_U0.stateTable2qpi_rsp_blk_n) begin
                            if (~stateTable2qpi_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.stateTable2qpi_rsp_U' written by process 'rocev2_top_rocev2_top.qp_interface_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.stateTable2qpi_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2qpi_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.stateTable2qpi_rsp_U' read by process 'rocev2_top_rocev2_top.qp_interface_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.stateTable2qpi_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                45 : begin
                    case(index2)
                    24: begin
                        if (~msn_table_0_U0.rxExh2msnTable_upd_req_blk_n) begin
                            if (~rxExh2msnTable_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rxExh2msnTable_upd_req_U' written by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rxExh2msnTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxExh2msnTable_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rxExh2msnTable_upd_req_U' read by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rxExh2msnTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~msn_table_0_U0.msnTable2rxExh_rsp_blk_n) begin
                            if (~msnTable2rxExh_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.msnTable2rxExh_rsp_U' written by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.msnTable2rxExh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~msnTable2rxExh_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.msnTable2rxExh_rsp_U' read by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.msnTable2rxExh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    36: begin
                        if (~msn_table_0_U0.txExh2msnTable_req_blk_n) begin
                            if (~txExh2msnTable_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.txExh2msnTable_req_U' written by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.txExh2msnTable_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txExh2msnTable_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.txExh2msnTable_req_U' read by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.txExh2msnTable_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~msn_table_0_U0.msnTable2txExh_rsp_blk_n) begin
                            if (~msnTable2txExh_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.msnTable2txExh_rsp_U' written by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.msnTable2txExh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~msnTable2txExh_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.msnTable2txExh_rsp_U' read by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.msnTable2txExh_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    17: begin
                        if (~msn_table_0_U0.if2msnTable_init_blk_n) begin
                            if (~if2msnTable_init_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.if2msnTable_init_U' written by process 'rocev2_top_rocev2_top.qp_interface_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.if2msnTable_init_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~if2msnTable_init_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.if2msnTable_init_U' read by process 'rocev2_top_rocev2_top.qp_interface_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.if2msnTable_init_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                46 : begin
                    case(index2)
                    39: begin
                        if (~merge_retrans_request_U0.tx2retrans_insertMeta_blk_n) begin
                            if (~tx2retrans_insertMeta_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx2retrans_insertMeta_U' written by process 'rocev2_top_rocev2_top.generate_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx2retrans_insertMeta_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx2retrans_insertMeta_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx2retrans_insertMeta_U' read by process 'rocev2_top_rocev2_top.generate_ibh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx2retrans_insertMeta_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    31: begin
                        if (~merge_retrans_request_U0.tx2retrans_insertAddrLen_blk_n) begin
                            if (~tx2retrans_insertAddrLen_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx2retrans_insertAddrLen_U' written by process 'rocev2_top_rocev2_top.local_req_handler_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx2retrans_insertAddrLen_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx2retrans_insertAddrLen_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx2retrans_insertAddrLen_U' read by process 'rocev2_top_rocev2_top.local_req_handler_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx2retrans_insertAddrLen_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    51: begin
                        if (~merge_retrans_request_U0.tx2retrans_insertRequest_blk_n) begin
                            if (~tx2retrans_insertRequest_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx2retrans_insertRequest_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx2retrans_insertRequest_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx2retrans_insertRequest_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx2retrans_insertRequest_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx2retrans_insertRequest_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                47 : begin
                    case(index2)
                    21: begin
                        if (~transport_timer_0_U0.rxClearTimer_req_blk_n) begin
                            if (~rxClearTimer_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rxClearTimer_req_U' written by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rxClearTimer_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxClearTimer_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rxClearTimer_req_U' read by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rxClearTimer_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    36: begin
                        if (~transport_timer_0_U0.txSetTimer_req_blk_n) begin
                            if (~txSetTimer_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.txSetTimer_req_U' written by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.txSetTimer_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txSetTimer_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.txSetTimer_req_U' read by process 'rocev2_top_rocev2_top.generate_exh_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.txSetTimer_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    51: begin
                        if (~transport_timer_0_U0.timer2retrans_req_blk_n) begin
                            if (~timer2retrans_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.timer2retrans_req_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.timer2retrans_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~timer2retrans_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.timer2retrans_req_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.timer2retrans_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                48 : begin
                    case(index2)
                    51: begin
                        if (~freelist_handler_0_U0.rt_releaseFifo_blk_n) begin
                            if (~rt_releaseFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_releaseFifo_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_releaseFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_releaseFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_releaseFifo_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_releaseFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~freelist_handler_0_U0.rt_freeListFifo_blk_n) begin
                            if (~rt_freeListFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_freeListFifo_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_freeListFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_freeListFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_freeListFifo_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_freeListFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                49 : begin
                    case(index2)
                    51: begin
                        if (~retrans_pointer_table_0_U0.rt_pointerUpdFifo_blk_n) begin
                            if (~rt_pointerUpdFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_pointerUpdFifo_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_pointerUpdFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_pointerUpdFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_pointerUpdFifo_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_pointerUpdFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~retrans_pointer_table_0_U0.rt_pointerReqFifo_blk_n) begin
                            if (~rt_pointerReqFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_pointerReqFifo_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_pointerReqFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_pointerReqFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_pointerReqFifo_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_pointerReqFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~retrans_pointer_table_0_U0.rt_pointerRspFifo_blk_n) begin
                            if (~rt_pointerRspFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_pointerRspFifo_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_pointerRspFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_pointerRspFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_pointerRspFifo_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_pointerRspFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                50 : begin
                    case(index2)
                    51: begin
                        if (~retrans_meta_table_0_U0.rt_metaReqFifo_blk_n) begin
                            if (~rt_metaReqFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_metaReqFifo_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_metaReqFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_metaReqFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_metaReqFifo_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_metaReqFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~retrans_meta_table_0_U0.rt_metaRspFifo_blk_n) begin
                            if (~rt_metaRspFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_metaRspFifo_U' written by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_metaRspFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_metaRspFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_metaRspFifo_U' read by process 'rocev2_top_rocev2_top.process_retransmissions_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_metaRspFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                51 : begin
                    case(index2)
                    21: begin
                        if (~process_retransmissions_0_U0.rx2retrans_upd_blk_n) begin
                            if (~rx2retrans_upd_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx2retrans_upd_U' written by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx2retrans_upd_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx2retrans_upd_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx2retrans_upd_U' read by process 'rocev2_top_rocev2_top.rx_ibh_fsm_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx2retrans_upd_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    49: begin
                        if (~process_retransmissions_0_U0.rt_pointerReqFifo_blk_n) begin
                            if (~rt_pointerReqFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_pointerReqFifo_U' written by process 'rocev2_top_rocev2_top.retrans_pointer_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_pointerReqFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_pointerReqFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_pointerReqFifo_U' read by process 'rocev2_top_rocev2_top.retrans_pointer_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_pointerReqFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~process_retransmissions_0_U0.rt_pointerRspFifo_blk_n) begin
                            if (~rt_pointerRspFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_pointerRspFifo_U' written by process 'rocev2_top_rocev2_top.retrans_pointer_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_pointerRspFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_pointerRspFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_pointerRspFifo_U' read by process 'rocev2_top_rocev2_top.retrans_pointer_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_pointerRspFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~process_retransmissions_0_U0.rt_pointerUpdFifo_blk_n) begin
                            if (~rt_pointerUpdFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_pointerUpdFifo_U' written by process 'rocev2_top_rocev2_top.retrans_pointer_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_pointerUpdFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_pointerUpdFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_pointerUpdFifo_U' read by process 'rocev2_top_rocev2_top.retrans_pointer_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_pointerUpdFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    24: begin
                        if (~process_retransmissions_0_U0.rx2retrans_req_blk_n) begin
                            if (~rx2retrans_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rx2retrans_req_U' written by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx2retrans_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx2retrans_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rx2retrans_req_U' read by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rx2retrans_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~process_retransmissions_0_U0.retrans2rx_init_blk_n) begin
                            if (~retrans2rx_init_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.retrans2rx_init_U' written by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.retrans2rx_init_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~retrans2rx_init_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.retrans2rx_init_U' read by process 'rocev2_top_rocev2_top.rx_exh_fsm_512_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.retrans2rx_init_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    47: begin
                        if (~process_retransmissions_0_U0.timer2retrans_req_blk_n) begin
                            if (~timer2retrans_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.timer2retrans_req_U' written by process 'rocev2_top_rocev2_top.transport_timer_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.timer2retrans_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~timer2retrans_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.timer2retrans_req_U' read by process 'rocev2_top_rocev2_top.transport_timer_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.timer2retrans_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    46: begin
                        if (~process_retransmissions_0_U0.tx2retrans_insertRequest_blk_n) begin
                            if (~tx2retrans_insertRequest_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.tx2retrans_insertRequest_U' written by process 'rocev2_top_rocev2_top.merge_retrans_request_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx2retrans_insertRequest_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tx2retrans_insertRequest_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.tx2retrans_insertRequest_U' read by process 'rocev2_top_rocev2_top.merge_retrans_request_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.tx2retrans_insertRequest_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    48: begin
                        if (~process_retransmissions_0_U0.rt_freeListFifo_blk_n) begin
                            if (~rt_freeListFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_freeListFifo_U' written by process 'rocev2_top_rocev2_top.freelist_handler_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_freeListFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_freeListFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_freeListFifo_U' read by process 'rocev2_top_rocev2_top.freelist_handler_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_freeListFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~process_retransmissions_0_U0.rt_releaseFifo_blk_n) begin
                            if (~rt_releaseFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_releaseFifo_U' written by process 'rocev2_top_rocev2_top.freelist_handler_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_releaseFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_releaseFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_releaseFifo_U' read by process 'rocev2_top_rocev2_top.freelist_handler_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_releaseFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    50: begin
                        if (~process_retransmissions_0_U0.rt_metaReqFifo_blk_n) begin
                            if (~rt_metaReqFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_metaReqFifo_U' written by process 'rocev2_top_rocev2_top.retrans_meta_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_metaReqFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_metaReqFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_metaReqFifo_U' read by process 'rocev2_top_rocev2_top.retrans_meta_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_metaReqFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~process_retransmissions_0_U0.rt_metaRspFifo_blk_n) begin
                            if (~rt_metaRspFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.rt_metaRspFifo_U' written by process 'rocev2_top_rocev2_top.retrans_meta_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_metaRspFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rt_metaRspFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.rt_metaRspFifo_U' read by process 'rocev2_top_rocev2_top.retrans_meta_table_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.rt_metaRspFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    31: begin
                        if (~process_retransmissions_0_U0.retransmitter2exh_eventFifo_blk_n) begin
                            if (~retransmitter2exh_eventFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'rocev2_top_rocev2_top.retransmitter2exh_eventFifo_U' written by process 'rocev2_top_rocev2_top.local_req_handler_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.retransmitter2exh_eventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~retransmitter2exh_eventFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'rocev2_top_rocev2_top.retransmitter2exh_eventFifo_U' read by process 'rocev2_top_rocev2_top.local_req_handler_0_U0'");
                                $fdisplay(fp, "Dependence_Channel_path rocev2_top_rocev2_top.retransmitter2exh_eventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        integer record_time;
        wait (dl_reset == 1);
        cycle_id = 1;
        record_time = 0;
        while (1) begin
            @ (negedge dl_clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                            record_time = $time;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end((cycle_id - 1),record_time);
                        @(negedge dl_clock);
                        @(negedge dl_clock);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
